module my_not (input in,
               output out);
   nand (out, in, in);
endmodule 
