module my_not (input in,
               output out);
   nand (out, in, 1);
endmodule 
