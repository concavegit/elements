module memory (input in, clock,
               output out);

   dff d0(in, clock, out);
endmodule
